library IEEE;
use IEEE.std_logic_1164.all;  
use IEEE.numeric_std.all;     

use work.pProc_bus_gb.all;
use work.pRegmap.all;

package pReg_ds_display_9 is

   -- range 0x00 .. 0x56
   --   (                                                    adr      upper    lower    size   default   accesstype)                                                     
   constant DISPCNT                        : regmap_type := (12#000#,  15,      0,        1,        0,   readwrite); -- LCD Control                                   2    R/W   
   constant DISPCNT_BG_Mode                : regmap_type := (12#000#,   2,      0,        1,        0,   readwrite); -- BG Mode                     (0-5=Video Mode 0-6, 7=Prohibited)
   constant DISPCNT_BG0_2D_3D              : regmap_type := (12#000#,   3,      3,        1,        0,   readwrite); -- A only BG0 2D/3D Selection (instead CGB Mode) (0=2D, 1=3D)
   constant DISPCNT_Tile_OBJ_Mapping       : regmap_type := (12#000#,   4,      4,        1,        0,   readwrite); -- Tile OBJ Mapping        (0=2D; max 32KB, 1=1D; max 32KB..256KB)
   constant DISPCNT_Bitmap_OBJ_2D_Dim      : regmap_type := (12#000#,   5,      5,        1,        0,   readwrite); -- Bitmap OBJ 2D-Dimension (0=128x512 dots, 1=256x256 dots)
   constant DISPCNT_Bitmap_OBJ_Mapping     : regmap_type := (12#000#,   6,      6,        1,        0,   readwrite); -- Bitmap OBJ Mapping      (0=2D; max 128KB, 1=1D; max 128KB..256KB)
   constant DISPCNT_Forced_Blank           : regmap_type := (12#000#,   7,      7,        1,        0,   readwrite); -- Forced Blank                (1=Allow FAST access to VRAM,Palette,OAM)
   constant DISPCNT_Screen_Display_BG0     : regmap_type := (12#000#,   8,      8,        1,        0,   readwrite); -- Screen Display BG0          (0=Off, 1=On)
   constant DISPCNT_Screen_Display_BG1     : regmap_type := (12#000#,   9,      9,        1,        0,   readwrite); -- Screen Display BG1          (0=Off, 1=On)
   constant DISPCNT_Screen_Display_BG2     : regmap_type := (12#000#,  10,     10,        1,        0,   readwrite); -- Screen Display BG2          (0=Off, 1=On)
   constant DISPCNT_Screen_Display_BG3     : regmap_type := (12#000#,  11,     11,        1,        0,   readwrite); -- Screen Display BG3          (0=Off, 1=On)
   constant DISPCNT_Screen_Display_OBJ     : regmap_type := (12#000#,  12,     12,        1,        0,   readwrite); -- Screen Display OBJ          (0=Off, 1=On)
   constant DISPCNT_Window_0_Display_Flag  : regmap_type := (12#000#,  13,     13,        1,        0,   readwrite); -- Window 0 Display Flag       (0=Off, 1=On)
   constant DISPCNT_Window_1_Display_Flag  : regmap_type := (12#000#,  14,     14,        1,        0,   readwrite); -- Window 1 Display Flag       (0=Off, 1=On)
   constant DISPCNT_OBJ_Wnd_Display_Flag   : regmap_type := (12#000#,  15,     15,        1,        0,   readwrite); -- OBJ Window Display Flag     (0=Off, 1=On)                                       
   constant DISPCNT_Display_Mode           : regmap_type := (12#000#,  17,     16,        1,        0,   readwrite); -- 16-17 A+B   Display Mode (Engine A: 0..3, Engine B: 0..1, GBA: Green Swap)
   constant DISPCNT_VRAM_block             : regmap_type := (12#000#,  19,     18,        1,        0,   readwrite); -- 18-19 A     VRAM block (0..3=VRAM A..D) (For Capture & above Display Mode=2)
   constant DISPCNT_Tile_OBJ_1D_Boundary   : regmap_type := (12#000#,  21,     20,        1,        0,   readwrite); -- 20-21 A+B   Tile OBJ 1D-Boundary   (see Bit4)
   constant DISPCNT_Bitmap_OBJ_1D_Boundary : regmap_type := (12#000#,  22,     22,        1,        0,   readwrite); -- 22    A     Bitmap OBJ 1D-Boundary (see Bit5-6)
   constant DISPCNT_OBJ_Process_H_Blank    : regmap_type := (12#000#,  23,     23,        1,        0,   readwrite); -- 23    A+B   OBJ Processing during H-Blank (was located in Bit5 on GBA)
   constant DISPCNT_Character_Base         : regmap_type := (12#000#,  26,     24,        1,        0,   readwrite); -- 24-26 A     Character Base (in 64K steps) (merged with 16K step in BGxCNT)
   constant DISPCNT_Screen_Base            : regmap_type := (12#000#,  29,     27,        1,        0,   readwrite); -- 27-29 A     Screen Base (in 64K steps) (merged with 2K step in BGxCNT)
   constant DISPCNT_BG_Extended_Palettes   : regmap_type := (12#000#,  30,     30,        1,        0,   readwrite); -- 30    A+B   BG Extended Palettes   (0=Disable, 1=Enable)
   constant DISPCNT_OBJ_Extended_Palettes  : regmap_type := (12#000#,  31,     31,        1,        0,   readwrite); -- 31    A+B   OBJ Extended Palettes  (0=Disable, 1=Enable
   
   constant DISPSTAT                       : regmap_type := (12#004#,  15,      0,        1, 16#0004#,   readwrite); -- General LCD Status (STAT,LYC)                 2    R/W
   constant DISPSTAT_V_Blank_flag          : regmap_type := (12#004#,   0,      0,        1,        0,   readonly ); -- V-Blank flag   (Read only) (1=VBlank) (set in line 160..226; not 227)
   constant DISPSTAT_H_Blank_flag          : regmap_type := (12#004#,   1,      1,        1,        0,   readonly ); -- H-Blank flag   (Read only) (1=HBlank) (toggled in all lines, 0..227)
   constant DISPSTAT_V_Counter_flag        : regmap_type := (12#004#,   2,      2,        1,        0,   readonly ); -- V-Counter flag (Read only) (1=Match)  (set in selected line)     (R)
   constant DISPSTAT_V_Blank_IRQ_Enable    : regmap_type := (12#004#,   3,      3,        1,        0,   readwrite); -- V-Blank IRQ Enable         (1=Enable)                          (R/W)
   constant DISPSTAT_H_Blank_IRQ_Enable    : regmap_type := (12#004#,   4,      4,        1,        0,   readwrite); -- H-Blank IRQ Enable         (1=Enable)                          (R/W)
   constant DISPSTAT_V_Counter_IRQ_Enable  : regmap_type := (12#004#,   5,      5,        1,        0,   readwrite); -- V-Counter IRQ Enable       (1=Enable)                          (R/W)
                                                                                                                     -- Not used (0) / DSi: LCD Initialization Ready (0=Busy, 1=Ready)   (R)
   constant DISPSTAT_V_Count_Setting8      : regmap_type := (12#004#,   7,      7,        1,        0,   readwrite); -- NDS: MSB of V-Vcount Setting (LYC.Bit8) (0..262)(R/W)
   constant DISPSTAT_V_Count_Setting       : regmap_type := (12#004#,  15,      8,        1,        0,   readwrite); -- V-Count Setting (LYC)      (0..227)                            (R/W)
                                           
   constant VCOUNT                         : regmap_type := (12#004#,  31,     16,        1,        0,   readwrite); -- Vertical Counter (LY)                         2    R  
                                           
   constant BG0CNT                         : regmap_type := (12#008#,  15,      0,        1,        0,   writeonly); -- BG0 Control                                   2    R/W
   constant BG0CNT_BG_Priority             : regmap_type := (12#008#,   1,      0,        1,        0,   readwrite); -- BG Priority           (0-3, 0=Highest)
   constant BG0CNT_Character_Base_Block    : regmap_type := (12#008#,   3,      2,        1,        0,   readwrite); -- Character Base Block  (0-3, in units of 16 KBytes) (=BG Tile Data)
   constant BG0CNT_UNUSED_4_5              : regmap_type := (12#008#,   5,      4,        1,        0,   readwrite); -- 4-5   Not used (must be zero)
   constant BG0CNT_Mosaic                  : regmap_type := (12#008#,   6,      6,        1,        0,   readwrite); -- Mosaic                (0=Disable, 1=Enable)
   constant BG0CNT_Colors_Palettes         : regmap_type := (12#008#,   7,      7,        1,        0,   readwrite); -- Colors/Palettes       (0=16/16, 1=256/1)
   constant BG0CNT_Screen_Base_Block       : regmap_type := (12#008#,  12,      8,        1,        0,   readwrite); -- Screen Base Block     (0-31, in units of 2 KBytes) (=BG Map Data)
   constant BG0CNT_Screen_Size             : regmap_type := (12#008#,  15,     14,        1,        0,   readwrite); -- Screen Size (0-3)
                                           
   constant BG1CNT                         : regmap_type := (12#00A#,  15,      0,        1,        0,   writeonly); -- BG1 Control                                   2    R/W
   constant BG1CNT_BG_Priority             : regmap_type := (12#00A#,   1,      0,        1,        0,   readwrite); -- BG Priority           (0-3, 0=Highest)
   constant BG1CNT_Character_Base_Block    : regmap_type := (12#00A#,   3,      2,        1,        0,   readwrite); -- Character Base Block  (0-3, in units of 16 KBytes) (=BG Tile Data)
   constant BG1CNT_UNUSED_4_5              : regmap_type := (12#00A#,   5,      4,        1,        0,   readwrite); -- 4-5   Not used (must be zero)
   constant BG1CNT_Mosaic                  : regmap_type := (12#00A#,   6,      6,        1,        0,   readwrite); -- Mosaic                (0=Disable, 1=Enable)
   constant BG1CNT_Colors_Palettes         : regmap_type := (12#00A#,   7,      7,        1,        0,   readwrite); -- Colors/Palettes       (0=16/16, 1=256/1)
   constant BG1CNT_Screen_Base_Block       : regmap_type := (12#00A#,  12,      8,        1,        0,   readwrite); -- Screen Base Block     (0-31, in units of 2 KBytes) (=BG Map Data)
   constant BG1CNT_Screen_Size             : regmap_type := (12#00A#,  15,     14,        1,        0,   readwrite); -- Screen Size (0-3)
                                           
   constant BG2CNT                         : regmap_type := (12#00C#,  15,      0,        1,        0,   readwrite); -- BG2 Control                                   2    R/W
   constant BG2CNT_BG_Priority             : regmap_type := (12#00C#,   1,      0,        1,        0,   readwrite); -- BG Priority           (0-3, 0=Highest)
   constant BG2CNT_Character_Base_Block    : regmap_type := (12#00C#,   3,      2,        1,        0,   readwrite); -- Character Base Block  (0-3, in units of 16 KBytes) (=BG Tile Data)
   constant BG2CNT_Mosaic                  : regmap_type := (12#00C#,   6,      6,        1,        0,   readwrite); -- Mosaic                (0=Disable, 1=Enable)
   constant BG2CNT_Colors_Palettes         : regmap_type := (12#00C#,   7,      7,        1,        0,   readwrite); -- Colors/Palettes       (0=16/16, 1=256/1)
   constant BG2CNT_Screen_Base_Block       : regmap_type := (12#00C#,  12,      8,        1,        0,   readwrite); -- Screen Base Block     (0-31, in units of 2 KBytes) (=BG Map Data)
   constant BG2CNT_Display_Area_Overflow   : regmap_type := (12#00C#,  13,     13,        1,        0,   readwrite); -- Display Area Overflow (0=Transparent, 1=Wraparound; BG2CNT/BG3CNT only)
   constant BG2CNT_Screen_Size             : regmap_type := (12#00C#,  15,     14,        1,        0,   readwrite); -- Screen Size (0-3)
                                           
   constant BG3CNT                         : regmap_type := (12#00E#,  15,      0,        1,        0,   readwrite); -- BG3 Control                                   2    R/W
   constant BG3CNT_BG_Priority             : regmap_type := (12#00E#,   1,      0,        1,        0,   readwrite); -- BG Priority           (0-3, 0=Highest)
   constant BG3CNT_Character_Base_Block    : regmap_type := (12#00E#,   3,      2,        1,        0,   readwrite); -- Character Base Block  (0-3, in units of 16 KBytes) (=BG Tile Data)
   constant BG3CNT_Mosaic                  : regmap_type := (12#00E#,   6,      6,        1,        0,   readwrite); -- Mosaic                (0=Disable, 1=Enable)
   constant BG3CNT_Colors_Palettes         : regmap_type := (12#00E#,   7,      7,        1,        0,   readwrite); -- Colors/Palettes       (0=16/16, 1=256/1)
   constant BG3CNT_Screen_Base_Block       : regmap_type := (12#00E#,  12,      8,        1,        0,   readwrite); -- Screen Base Block     (0-31, in units of 2 KBytes) (=BG Map Data)
   constant BG3CNT_Display_Area_Overflow   : regmap_type := (12#00E#,  13,     13,        1,        0,   readwrite); -- Display Area Overflow (0=Transparent, 1=Wraparound; BG2CNT/BG3CNT only)
   constant BG3CNT_Screen_Size             : regmap_type := (12#00E#,  15,     14,        1,        0,   readwrite); -- Screen Size (0-3)
                                           
   constant BG0HOFS                        : regmap_type := (12#010#,  15,      0,        1,        0,   writeonly); -- BG0 X-Offset                                  2    W  
   constant BG0VOFS                        : regmap_type := (12#012#,  15,      0,        1,        0,   writeonly); -- BG0 Y-Offset                                  2    W  
   constant BG1HOFS                        : regmap_type := (12#014#,  15,      0,        1,        0,   writeonly); -- BG1 X-Offset                                  2    W  
   constant BG1VOFS                        : regmap_type := (12#016#,  15,      0,        1,        0,   writeonly); -- BG1 Y-Offset                                  2    W  
   constant BG2HOFS                        : regmap_type := (12#018#,  15,      0,        1,        0,   writeonly); -- BG2 X-Offset                                  2    W  
   constant BG2VOFS                        : regmap_type := (12#01A#,  15,      0,        1,        0,   writeonly); -- BG2 Y-Offset                                  2    W  
   constant BG3HOFS                        : regmap_type := (12#01C#,  15,      0,        1,        0,   writeonly); -- BG3 X-Offset                                  2    W  
   constant BG3VOFS                        : regmap_type := (12#01E#,  15,      0,        1,        0,   writeonly); -- BG3 Y-Offset                                  2    W  
                                           
   constant BG2RotScaleParDX               : regmap_type := (12#020#,  15,      0,        1,      256,   writeonly); -- BG2 Rotation/Scaling Parameter A (dx)         2    W  
   constant BG2RotScaleParDMX              : regmap_type := (12#020#,  31,     16,        1,        0,   writeonly); -- BG2 Rotation/Scaling Parameter B (dmx)        2    W  
   constant BG2RotScaleParDY               : regmap_type := (12#024#,  15,      0,        1,        0,   writeonly); -- BG2 Rotation/Scaling Parameter C (dy)         2    W  
   constant BG2RotScaleParDMY              : regmap_type := (12#024#,  31,     16,        1,      256,   writeonly); -- BG2 Rotation/Scaling Parameter D (dmy)        2    W  
   constant BG2RefX                        : regmap_type := (12#028#,  27,      0,        1,        0,   writeonly); -- BG2 Reference Point X-Coordinate              4    W  
   constant BG2RefY                        : regmap_type := (12#02C#,  27,      0,        1,        0,   writeonly); -- BG2 Reference Point Y-Coordinate              4    W  
                                           
   constant BG3RotScaleParDX               : regmap_type := (12#030#,  15,      0,        1,      256,   writeonly); -- BG3 Rotation/Scaling Parameter A (dx)         2    W  
   constant BG3RotScaleParDMX              : regmap_type := (12#030#,  31,     16,        1,        0,   writeonly); -- BG3 Rotation/Scaling Parameter B (dmx)        2    W  
   constant BG3RotScaleParDY               : regmap_type := (12#034#,  15,      0,        1,        0,   writeonly); -- BG3 Rotation/Scaling Parameter C (dy)         2    W  
   constant BG3RotScaleParDMY              : regmap_type := (12#034#,  31,     16,        1,      256,   writeonly); -- BG3 Rotation/Scaling Parameter D (dmy)        2    W  
   constant BG3RefX                        : regmap_type := (12#038#,  27,      0,        1,        0,   writeonly); -- BG3 Reference Point X-Coordinate              4    W  
   constant BG3RefY                        : regmap_type := (12#03C#,  27,      0,        1,        0,   writeonly); -- BG3 Reference Point Y-Coordinate              4    W  
                                           
   constant WIN0H                          : regmap_type := (12#040#,  15,      0,        1,        0,   writeonly); -- Window 0 Horizontal Dimensions                2    W  
   constant WIN0H_X2                       : regmap_type := (12#040#,   7,      0,        1,        0,   writeonly); -- Window 0 Horizontal Dimensions                2    W  
   constant WIN0H_X1                       : regmap_type := (12#040#,  15,      8,        1,        0,   writeonly); -- Window 0 Horizontal Dimensions                2    W  
                                           
   constant WIN1H                          : regmap_type := (12#040#,  31,     16,        1,        0,   writeonly); -- Window 1 Horizontal Dimensions                2    W  
   constant WIN1H_X2                       : regmap_type := (12#040#,  23,     16,        1,        0,   writeonly); -- Window 1 Horizontal Dimensions                2    W  
   constant WIN1H_X1                       : regmap_type := (12#040#,  31,     24,        1,        0,   writeonly); -- Window 1 Horizontal Dimensions                2    W  
                                           
   constant WIN0V                          : regmap_type := (12#044#,  15,      0,        1,        0,   writeonly); -- Window 0 Vertical Dimensions                  2    W  
   constant WIN0V_Y2                       : regmap_type := (12#044#,   7,      0,        1,        0,   writeonly); -- Window 0 Vertical Dimensions                  2    W  
   constant WIN0V_Y1                       : regmap_type := (12#044#,  15,      8,        1,        0,   writeonly); -- Window 0 Vertical Dimensions                  2    W  
                                                                       
   constant WIN1V                          : regmap_type := (12#044#,  31,     16,        1,        0,   writeonly); -- Window 1 Vertical Dimensions                  2    W  
   constant WIN1V_Y2                       : regmap_type := (12#044#,  23,     16,        1,        0,   writeonly); -- Window 1 Vertical Dimensions                  2    W  
   constant WIN1V_Y1                       : regmap_type := (12#044#,  31,     24,        1,        0,   writeonly); -- Window 1 Vertical Dimensions                  2    W  
                                           
   constant WININ                          : regmap_type := (12#048#,  15,      0,        1,        0,   writeonly); -- Inside of Window 0 and 1                      2    R/W
   constant WININ_Window_0_BG0_Enable      : regmap_type := (12#048#,   0,      0,        1,        0,   readwrite); -- 0-3   Window_0_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_0_BG1_Enable      : regmap_type := (12#048#,   1,      1,        1,        0,   readwrite); -- 0-3   Window_0_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_0_BG2_Enable      : regmap_type := (12#048#,   2,      2,        1,        0,   readwrite); -- 0-3   Window_0_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_0_BG3_Enable      : regmap_type := (12#048#,   3,      3,        1,        0,   readwrite); -- 0-3   Window_0_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_0_OBJ_Enable      : regmap_type := (12#048#,   4,      4,        1,        0,   readwrite); -- 4     Window_0_OBJ_Enable         (0=No Display, 1=Display)
   constant WININ_Window_0_Special_Effect  : regmap_type := (12#048#,   5,      5,        1,        0,   readwrite); -- 5     Window_0_Special_Effect     (0=Disable, 1=Enable)
   constant WININ_Window_1_BG0_Enable      : regmap_type := (12#048#,   8,      8,        1,        0,   readwrite); -- 8-11  Window_1_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_1_BG1_Enable      : regmap_type := (12#048#,   9,      9,        1,        0,   readwrite); -- 8-11  Window_1_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_1_BG2_Enable      : regmap_type := (12#048#,  10,     10,        1,        0,   readwrite); -- 8-11  Window_1_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_1_BG3_Enable      : regmap_type := (12#048#,  11,     11,        1,        0,   readwrite); -- 8-11  Window_1_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WININ_Window_1_OBJ_Enable      : regmap_type := (12#048#,  12,     12,        1,        0,   readwrite); -- 12    Window_1_OBJ_Enable         (0=No Display, 1=Display)
   constant WININ_Window_1_Special_Effect  : regmap_type := (12#048#,  13,     13,        1,        0,   readwrite); -- 13    Window_1_Special_Effect     (0=Disable, 1=Enable)
                                           
   constant WINOUT                         : regmap_type := (12#048#,  31,     16,        1,        0,   writeonly); -- Inside of OBJ Window & Outside of Windows     2    R/W
   constant WINOUT_Outside_BG0_Enable      : regmap_type := (12#048#,  16,     16,        1,        0,   readwrite); -- 0-3   Outside_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Outside_BG1_Enable      : regmap_type := (12#048#,  17,     17,        1,        0,   readwrite); -- 0-3   Outside_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Outside_BG2_Enable      : regmap_type := (12#048#,  18,     18,        1,        0,   readwrite); -- 0-3   Outside_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Outside_BG3_Enable      : regmap_type := (12#048#,  19,     19,        1,        0,   readwrite); -- 0-3   Outside_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Outside_OBJ_Enable      : regmap_type := (12#048#,  20,     20,        1,        0,   readwrite); -- 4     Outside_OBJ_Enable         (0=No Display, 1=Display)
   constant WINOUT_Outside_Special_Effect  : regmap_type := (12#048#,  21,     21,        1,        0,   readwrite); -- 5     Outside_Special_Effect     (0=Disable, 1=Enable)
   constant WINOUT_Objwnd_BG0_Enable       : regmap_type := (12#048#,  24,     24,        1,        0,   readwrite); -- 8-11  object window_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Objwnd_BG1_Enable       : regmap_type := (12#048#,  25,     25,        1,        0,   readwrite); -- 8-11  object window_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Objwnd_BG2_Enable       : regmap_type := (12#048#,  26,     26,        1,        0,   readwrite); -- 8-11  object window_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Objwnd_BG3_Enable       : regmap_type := (12#048#,  27,     27,        1,        0,   readwrite); -- 8-11  object window_BG0_BG3_Enable     (0=No Display, 1=Display)
   constant WINOUT_Objwnd_OBJ_Enable       : regmap_type := (12#048#,  28,     28,        1,        0,   readwrite); -- 12    object window_OBJ_Enable         (0=No Display, 1=Display)
   constant WINOUT_Objwnd_Special_Effect   : regmap_type := (12#048#,  29,     29,        1,        0,   readwrite); -- 13    object window_Special_Effect     (0=Disable, 1=Enable)
                                           
   constant MOSAIC                         : regmap_type := (12#04C#,  15,      0,        1,        0,   writeonly); -- Mosaic Size                                   2    W  
   constant MOSAIC_BG_Mosaic_H_Size        : regmap_type := (12#04C#,   3,      0,        1,        0,   writeonly); --   0-3   BG_Mosaic_H_Size  (minus 1)  
   constant MOSAIC_BG_Mosaic_V_Size        : regmap_type := (12#04C#,   7,      4,        1,        0,   writeonly); --   4-7   BG_Mosaic_V_Size  (minus 1)  
   constant MOSAIC_OBJ_Mosaic_H_Size       : regmap_type := (12#04C#,  11,      8,        1,        0,   writeonly); --   8-11  OBJ_Mosaic_H_Size (minus 1)  
   constant MOSAIC_OBJ_Mosaic_V_Size       : regmap_type := (12#04C#,  15,     12,        1,        0,   writeonly); --   12-15 OBJ_Mosaic_V_Size (minus 1)  
                                           
   constant BLDCNT                         : regmap_type := (12#050#,  13,      0,        1,        0,   readwrite); -- Color Special Effects Selection               2    R/W
   constant BLDCNT_BG0_1st_Target_Pixel    : regmap_type := (12#050#,   0,      0,        1,        0,   readwrite); -- 0      (Background 0)
   constant BLDCNT_BG1_1st_Target_Pixel    : regmap_type := (12#050#,   1,      1,        1,        0,   readwrite); -- 1      (Background 1)
   constant BLDCNT_BG2_1st_Target_Pixel    : regmap_type := (12#050#,   2,      2,        1,        0,   readwrite); -- 2      (Background 2)
   constant BLDCNT_BG3_1st_Target_Pixel    : regmap_type := (12#050#,   3,      3,        1,        0,   readwrite); -- 3      (Background 3)
   constant BLDCNT_OBJ_1st_Target_Pixel    : regmap_type := (12#050#,   4,      4,        1,        0,   readwrite); -- 4      (Top-most OBJ pixel)
   constant BLDCNT_BD_1st_Target_Pixel     : regmap_type := (12#050#,   5,      5,        1,        0,   readwrite); -- 5      (Backdrop)
   constant BLDCNT_Color_Special_Effect    : regmap_type := (12#050#,   7,      6,        1,        0,   readwrite); -- 6-7    (0-3, see below) 0 = None (Special effects disabled), 1 = Alpha Blending (1st+2nd Target mixed), 2 = Brightness Increase (1st Target becomes whiter), 3 = Brightness Decrease (1st Target becomes blacker)
   constant BLDCNT_BG0_2nd_Target_Pixel    : regmap_type := (12#050#,   8,      8,        1,        0,   readwrite); -- 8      (Background 0)
   constant BLDCNT_BG1_2nd_Target_Pixel    : regmap_type := (12#050#,   9,      9,        1,        0,   readwrite); -- 9      (Background 1)
   constant BLDCNT_BG2_2nd_Target_Pixel    : regmap_type := (12#050#,  10,     10,        1,        0,   readwrite); -- 10     (Background 2)
   constant BLDCNT_BG3_2nd_Target_Pixel    : regmap_type := (12#050#,  11,     11,        1,        0,   readwrite); -- 11     (Background 3)
   constant BLDCNT_OBJ_2nd_Target_Pixel    : regmap_type := (12#050#,  12,     12,        1,        0,   readwrite); -- 12     (Top-most OBJ pixel)
   constant BLDCNT_BD_2nd_Target_Pixel     : regmap_type := (12#050#,  13,     13,        1,        0,   readwrite); -- 13     (Backdrop)
                                           
   constant BLDALPHA                       : regmap_type := (12#050#,  28,     16,        1,        0,   writeonly); -- Alpha Blending Coefficients                   2    W  
   constant BLDALPHA_EVA_Coefficient       : regmap_type := (12#050#,  20,     16,        1,        0,   readwrite); -- 0-4   (1st Target) (0..16 = 0/16..16/16, 17..31=16/16)
   constant BLDALPHA_EVB_Coefficient       : regmap_type := (12#050#,  28,     24,        1,        0,   readwrite); -- 8-12  (2nd Target) (0..16 = 0/16..16/16, 17..31=16/16)
                                           
   constant BLDY                           : regmap_type := (12#054#,   4,      0,        1,        0,   writeonly); -- Brightness (Fade-In/Out) Coefficient  0-4   EVY Coefficient (Brightness) (0..16 = 0/16..16/16, 17..31=16/16 
                                           
   constant DISPCAPCNT                     : regmap_type := (12#064#,  31,      0,        1,        0,   writeonly); -- Alpha Blending Coefficients                   2    W  
   constant DISPCAPCNT_EVA                 : regmap_type := (12#064#,   4,      0,        1,        0,   writeonly); -- 0-4   EVA               (0..16 = Blending Factor for Source A)
   constant DISPCAPCNT_EVB                 : regmap_type := (12#064#,  12,      8,        1,        0,   writeonly); -- 8-12  EVB               (0..16 = Blending Factor for Source B)
   constant DISPCAPCNT_VRAM_Write_Block    : regmap_type := (12#064#,  17,     16,        1,        0,   writeonly); -- 16-17 VRAM Write Block  (0..3 = VRAM A..D) (VRAM must be allocated to LCDC)
   constant DISPCAPCNT_VRAM_Write_Offset   : regmap_type := (12#064#,  19,     18,        1,        0,   writeonly); -- 18-19 VRAM Write Offset (0=00000h, 0=08000h, 0=10000h, 0=18000h)
   constant DISPCAPCNT_Capture_Size        : regmap_type := (12#064#,  21,     20,        1,        0,   writeonly); -- 20-21 Capture Size      (0=128x128, 1=256x64, 2=256x128, 3=256x192 dots)
   constant DISPCAPCNT_Source_A            : regmap_type := (12#064#,  24,     24,        1,        0,   writeonly); -- 24    Source A          (0=Graphics Screen BG+3D+OBJ, 1=3D Screen)
   constant DISPCAPCNT_Source_B            : regmap_type := (12#064#,  25,     25,        1,        0,   writeonly); -- 25    Source B          (0=VRAM, 1=Main Memory Display FIFO)
   constant DISPCAPCNT_VRAM_Read_Offset    : regmap_type := (12#064#,  27,     26,        1,        0,   writeonly); -- 26-27 VRAM Read Offset  (0=00000h, 0=08000h, 0=10000h, 0=18000h)
   constant DISPCAPCNT_Capture_Source      : regmap_type := (12#064#,  30,     29,        1,        0,   writeonly); -- 29-30 Capture Source    (0=Source A, 1=Source B, 2/3=Sources A+B blended)
   constant DISPCAPCNT_Capture_Enable      : regmap_type := (12#064#,  31,     31,        1,        0,   writeonly); -- 31    Capture Enable    (0=Disable/Ready, 1=Enable/Busy)
                                           
   constant DISP_MMEM_FIFO                 : regmap_type := (12#068#,  31,      0,        1,        0,   writeonly); -- Main Memory Display FIFO (R?/W)
                                           
   constant MASTER_BRIGHT                  : regmap_type := (12#06C#,  15,      0,        1,        0,   writeonly); -- Alpha Blending Coefficients                   2    W  
   constant MASTER_BRIGHT_Factor           : regmap_type := (12#06C#,   4,      0,        1,        0,   writeonly); -- Factor used for 6bit R,G,B Intensities (0-16, values >16 same as 16)
   constant MASTER_BRIGHT_Mode             : regmap_type := (12#06C#,  15,     14,        1,        0,   writeonly); -- Mode (0=Disable, 1=Up, 2=Down, 3=Reserved)
 
  
   
end package;

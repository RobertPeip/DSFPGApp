library IEEE;
use IEEE.std_logic_1164.all;  
use IEEE.numeric_std.all;     

use work.pProc_bus_gb.all;
use work.pRegmap.all;

package pReg_ds_sound_7 is

   -- range 0x400 .. 0x51F
   --   (                                                              adr      upper    lower    size   default   accesstype)                                     
   constant SOUND0CNT                                : regmap_type := (16#400#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND0CNT_Volume_Mul                     : regmap_type := (16#400#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND0CNT_Volume_Div                     : regmap_type := (16#400#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND0CNT_Hold                           : regmap_type := (16#400#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND0CNT_Panning                        : regmap_type := (16#400#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND0CNT_Wave_Duty                      : regmap_type := (16#400#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND0CNT_Repeat_Mode                    : regmap_type := (16#400#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND0CNT_Format                         : regmap_type := (16#400#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND0CNT_Start_Status                   : regmap_type := (16#400#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND0SAD                                : regmap_type := (16#404#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND0TMR                                : regmap_type := (16#408#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND0PNT                                : regmap_type := (16#408#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND0LEN                                : regmap_type := (16#40C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
  
   constant SOUND1CNT                                : regmap_type := (16#410#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND1CNT_Volume_Mul                     : regmap_type := (16#410#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND1CNT_Volume_Div                     : regmap_type := (16#410#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND1CNT_Hold                           : regmap_type := (16#410#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND1CNT_Panning                        : regmap_type := (16#410#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND1CNT_Wave_Duty                      : regmap_type := (16#410#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND1CNT_Repeat_Mode                    : regmap_type := (16#410#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND1CNT_Format                         : regmap_type := (16#410#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND1CNT_Start_Status                   : regmap_type := (16#410#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND1SAD                                : regmap_type := (16#414#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND1TMR                                : regmap_type := (16#418#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND1PNT                                : regmap_type := (16#418#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND1LEN                                : regmap_type := (16#41C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND2CNT                                : regmap_type := (16#420#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND2CNT_Volume_Mul                     : regmap_type := (16#420#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND2CNT_Volume_Div                     : regmap_type := (16#420#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND2CNT_Hold                           : regmap_type := (16#420#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND2CNT_Panning                        : regmap_type := (16#420#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND2CNT_Wave_Duty                      : regmap_type := (16#420#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND2CNT_Repeat_Mode                    : regmap_type := (16#420#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND2CNT_Format                         : regmap_type := (16#420#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND2CNT_Start_Status                   : regmap_type := (16#420#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND2SAD                                : regmap_type := (16#424#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND2TMR                                : regmap_type := (16#428#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND2PNT                                : regmap_type := (16#428#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND2LEN                                : regmap_type := (16#42C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND3CNT                                : regmap_type := (16#430#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND3CNT_Volume_Mul                     : regmap_type := (16#430#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND3CNT_Volume_Div                     : regmap_type := (16#430#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND3CNT_Hold                           : regmap_type := (16#430#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND3CNT_Panning                        : regmap_type := (16#430#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND3CNT_Wave_Duty                      : regmap_type := (16#430#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND3CNT_Repeat_Mode                    : regmap_type := (16#430#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND3CNT_Format                         : regmap_type := (16#430#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND3CNT_Start_Status                   : regmap_type := (16#430#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND3SAD                                : regmap_type := (16#434#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND3TMR                                : regmap_type := (16#438#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND3PNT                                : regmap_type := (16#438#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND3LEN                                : regmap_type := (16#43C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND4CNT                                : regmap_type := (16#440#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND4CNT_Volume_Mul                     : regmap_type := (16#440#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND4CNT_Volume_Div                     : regmap_type := (16#440#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND4CNT_Hold                           : regmap_type := (16#440#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND4CNT_Panning                        : regmap_type := (16#440#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND4CNT_Wave_Duty                      : regmap_type := (16#440#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND4CNT_Repeat_Mode                    : regmap_type := (16#440#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND4CNT_Format                         : regmap_type := (16#440#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND4CNT_Start_Status                   : regmap_type := (16#440#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND4SAD                                : regmap_type := (16#444#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND4TMR                                : regmap_type := (16#448#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND4PNT                                : regmap_type := (16#448#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND4LEN                                : regmap_type := (16#44C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND5CNT                                : regmap_type := (16#450#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND5CNT_Volume_Mul                     : regmap_type := (16#450#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND5CNT_Volume_Div                     : regmap_type := (16#450#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND5CNT_Hold                           : regmap_type := (16#450#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND5CNT_Panning                        : regmap_type := (16#450#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND5CNT_Wave_Duty                      : regmap_type := (16#450#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND5CNT_Repeat_Mode                    : regmap_type := (16#450#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND5CNT_Format                         : regmap_type := (16#450#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND5CNT_Start_Status                   : regmap_type := (16#450#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND5SAD                                : regmap_type := (16#454#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND5TMR                                : regmap_type := (16#458#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND5PNT                                : regmap_type := (16#458#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND5LEN                                : regmap_type := (16#45C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND6CNT                                : regmap_type := (16#460#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND6CNT_Volume_Mul                     : regmap_type := (16#460#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND6CNT_Volume_Div                     : regmap_type := (16#460#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND6CNT_Hold                           : regmap_type := (16#460#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND6CNT_Panning                        : regmap_type := (16#460#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND6CNT_Wave_Duty                      : regmap_type := (16#460#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND6CNT_Repeat_Mode                    : regmap_type := (16#460#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND6CNT_Format                         : regmap_type := (16#460#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND6CNT_Start_Status                   : regmap_type := (16#460#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND6SAD                                : regmap_type := (16#464#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND6TMR                                : regmap_type := (16#468#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND6PNT                                : regmap_type := (16#468#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND6LEN                                : regmap_type := (16#46C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND7CNT                                : regmap_type := (16#470#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND7CNT_Volume_Mul                     : regmap_type := (16#470#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND7CNT_Volume_Div                     : regmap_type := (16#470#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND7CNT_Hold                           : regmap_type := (16#470#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND7CNT_Panning                        : regmap_type := (16#470#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND7CNT_Wave_Duty                      : regmap_type := (16#470#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND7CNT_Repeat_Mode                    : regmap_type := (16#470#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND7CNT_Format                         : regmap_type := (16#470#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND7CNT_Start_Status                   : regmap_type := (16#470#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND7SAD                                : regmap_type := (16#474#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND7TMR                                : regmap_type := (16#478#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND7PNT                                : regmap_type := (16#478#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND7LEN                                : regmap_type := (16#47C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND8CNT                                : regmap_type := (16#480#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND8CNT_Volume_Mul                     : regmap_type := (16#480#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND8CNT_Volume_Div                     : regmap_type := (16#480#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND8CNT_Hold                           : regmap_type := (16#480#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND8CNT_Panning                        : regmap_type := (16#480#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND8CNT_Wave_Duty                      : regmap_type := (16#480#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND8CNT_Repeat_Mode                    : regmap_type := (16#480#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND8CNT_Format                         : regmap_type := (16#480#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND8CNT_Start_Status                   : regmap_type := (16#480#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND8SAD                                : regmap_type := (16#484#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND8TMR                                : regmap_type := (16#488#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND8PNT                                : regmap_type := (16#488#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND8LEN                                : regmap_type := (16#48C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND9CNT                                : regmap_type := (16#490#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND9CNT_Volume_Mul                     : regmap_type := (16#490#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND9CNT_Volume_Div                     : regmap_type := (16#490#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND9CNT_Hold                           : regmap_type := (16#490#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND9CNT_Panning                        : regmap_type := (16#490#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND9CNT_Wave_Duty                      : regmap_type := (16#490#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND9CNT_Repeat_Mode                    : regmap_type := (16#490#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND9CNT_Format                         : regmap_type := (16#490#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND9CNT_Start_Status                   : regmap_type := (16#490#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND9SAD                                : regmap_type := (16#494#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND9TMR                                : regmap_type := (16#498#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND9PNT                                : regmap_type := (16#498#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND9LEN                                : regmap_type := (16#49C#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND10CNT                               : regmap_type := (16#4A0#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND10CNT_Volume_Mul                    : regmap_type := (16#4A0#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND10CNT_Volume_Div                    : regmap_type := (16#4A0#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND10CNT_Hold                          : regmap_type := (16#4A0#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND10CNT_Panning                       : regmap_type := (16#4A0#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND10CNT_Wave_Duty                     : regmap_type := (16#4A0#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND10CNT_Repeat_Mode                   : regmap_type := (16#4A0#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND10CNT_Format                        : regmap_type := (16#4A0#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND10CNT_Start_Status                  : regmap_type := (16#4A0#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND10SAD                               : regmap_type := (16#4A4#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND10TMR                               : regmap_type := (16#4A8#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND10PNT                               : regmap_type := (16#4A8#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND10LEN                               : regmap_type := (16#4AC#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND11CNT                               : regmap_type := (16#4B0#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND11CNT_Volume_Mul                    : regmap_type := (16#4B0#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND11CNT_Volume_Div                    : regmap_type := (16#4B0#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND11CNT_Hold                          : regmap_type := (16#4B0#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND11CNT_Panning                       : regmap_type := (16#4B0#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND11CNT_Wave_Duty                     : regmap_type := (16#4B0#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND11CNT_Repeat_Mode                   : regmap_type := (16#4B0#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND11CNT_Format                        : regmap_type := (16#4B0#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND11CNT_Start_Status                  : regmap_type := (16#4B0#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND11SAD                               : regmap_type := (16#4B4#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND11TMR                               : regmap_type := (16#4B8#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND11PNT                               : regmap_type := (16#4B8#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND11LEN                               : regmap_type := (16#4BC#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND12CNT                               : regmap_type := (16#4C0#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND12CNT_Volume_Mul                    : regmap_type := (16#4C0#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND12CNT_Volume_Div                    : regmap_type := (16#4C0#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND12CNT_Hold                          : regmap_type := (16#4C0#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND12CNT_Panning                       : regmap_type := (16#4C0#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND12CNT_Wave_Duty                     : regmap_type := (16#4C0#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND12CNT_Repeat_Mode                   : regmap_type := (16#4C0#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND12CNT_Format                        : regmap_type := (16#4C0#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND12CNT_Start_Status                  : regmap_type := (16#4C0#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND12SAD                               : regmap_type := (16#4C4#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND12TMR                               : regmap_type := (16#4C8#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND12PNT                               : regmap_type := (16#4C8#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND12LEN                               : regmap_type := (16#4CC#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND13CNT                               : regmap_type := (16#4D0#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND13CNT_Volume_Mul                    : regmap_type := (16#4D0#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND13CNT_Volume_Div                    : regmap_type := (16#4D0#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND13CNT_Hold                          : regmap_type := (16#4D0#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND13CNT_Panning                       : regmap_type := (16#4D0#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND13CNT_Wave_Duty                     : regmap_type := (16#4D0#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND13CNT_Repeat_Mode                   : regmap_type := (16#4D0#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND13CNT_Format                        : regmap_type := (16#4D0#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND13CNT_Start_Status                  : regmap_type := (16#4D0#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND13SAD                               : regmap_type := (16#4D4#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND13TMR                               : regmap_type := (16#4D8#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND13PNT                               : regmap_type := (16#4D8#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND13LEN                               : regmap_type := (16#4DC#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND14CNT                               : regmap_type := (16#4E0#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND14CNT_Volume_Mul                    : regmap_type := (16#4E0#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND14CNT_Volume_Div                    : regmap_type := (16#4E0#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND14CNT_Hold                          : regmap_type := (16#4E0#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND14CNT_Panning                       : regmap_type := (16#4E0#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND14CNT_Wave_Duty                     : regmap_type := (16#4E0#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND14CNT_Repeat_Mode                   : regmap_type := (16#4E0#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND14CNT_Format                        : regmap_type := (16#4E0#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND14CNT_Start_Status                  : regmap_type := (16#4E0#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND14SAD                               : regmap_type := (16#4E4#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND14TMR                               : regmap_type := (16#4E8#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND14PNT                               : regmap_type := (16#4E8#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND14LEN                               : regmap_type := (16#4EC#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUND15CNT                               : regmap_type := (16#4F0#,  31,      0,        1,        0,   writeonly); -- SOUNDxCNT - Sound Channel X Control Register (R/W)
   constant SOUND15CNT_Volume_Mul                    : regmap_type := (16#4F0#,   6,      0,        1,        0,   readwrite); -- 0-6    Volume Mul   (0..127=silent..loud)
   constant SOUND15CNT_Volume_Div                    : regmap_type := (16#4F0#,   9,      8,        1,        0,   readwrite); -- 8-9    Volume Div   (0=Normal, 1=Div2, 2=Div4, 3=Div16)
   constant SOUND15CNT_Hold                          : regmap_type := (16#4F0#,  15,     15,        1,        0,   readwrite); -- 15     Hold         (0=Normal, 1=Hold last sample after one-shot sound)
   constant SOUND15CNT_Panning                       : regmap_type := (16#4F0#,  22,     16,        1,        0,   readwrite); -- 16-22  Panning      (0..127=left..right) (64=half volume on both speakers)
   constant SOUND15CNT_Wave_Duty                     : regmap_type := (16#4F0#,  26,     24,        1,        0,   readwrite); -- 24-26  Wave Duty    (0..7) ;HIGH=(N+1)*12.5%, LOW=(7-N)*12.5% (PSG only)
   constant SOUND15CNT_Repeat_Mode                   : regmap_type := (16#4F0#,  28,     27,        1,        0,   readwrite); -- 27-28  Repeat Mode  (0=Manual, 1=Loop Infinite, 2=One-Shot, 3=Prohibited)
   constant SOUND15CNT_Format                        : regmap_type := (16#4F0#,  30,     29,        1,        0,   readwrite); -- 29-30  Format       (0=PCM8, 1=PCM16, 2=IMA-ADPCM, 3=PSG/Noise)
   constant SOUND15CNT_Start_Status                  : regmap_type := (16#4F0#,  31,     31,        1,        0,   readwrite); -- 31     Start/Status (0=Stop, 1=Start/Busy)
   constant SOUND15SAD                               : regmap_type := (16#4F4#,  26,      0,        1,        0,   writeonly); -- SOUNDxSAD - Sound Channel X Data Source Register (W)
   constant SOUND15TMR                               : regmap_type := (16#4F8#,  15,      0,        1,        0,   writeonly); -- SOUNDxTMR - Sound Channel X Timer Register (W)
   constant SOUND15PNT                               : regmap_type := (16#4F8#,  31,     16,        1,        0,   writeonly); -- SOUNDxPNT - Sound Channel X Loopstart Register (W)
   constant SOUND15LEN                               : regmap_type := (16#4FC#,  21,     16,        1,        0,   writeonly); -- SOUNDxLEN - Sound Channel X Length Register (W)
   
   constant SOUNDCNT                                 : regmap_type := (16#500#,  15,      0,        1,        0,   writeonly); -- 
   constant SOUNDCNT_Master_Volume                   : regmap_type := (16#500#,   6,      0,        1,        0,   readwrite); -- Bit0-6   Master Volume       (0..127=silent..loud)
   constant SOUNDCNT_Left_Output_from                : regmap_type := (16#500#,   9,      8,        1,        0,   readwrite); -- Bit8-9   Left Output from    (0=Left Mixer, 1=Ch1, 2=Ch3, 3=Ch1+Ch3)
   constant SOUNDCNT_Right_Output_from               : regmap_type := (16#500#,  11,     10,        1,        0,   readwrite); -- Bit10-11 Right Output from   (0=Right Mixer, 1=Ch1, 2=Ch3, 3=Ch1+Ch3)
   constant SOUNDCNT_Output_Ch1_to_Mixer             : regmap_type := (16#500#,  12,     12,        1,        0,   readwrite); -- Bit12    Output Ch1 to Mixer (0=Yes, 1=No) (both Left/Right)
   constant SOUNDCNT_Output_Ch3_to_Mixer             : regmap_type := (16#500#,  13,     13,        1,        0,   readwrite); -- Bit13    Output Ch3 to Mixer (0=Yes, 1=No) (both Left/Right)
   constant SOUNDCNT_Master_Enable                   : regmap_type := (16#500#,  15,     15,        1,        0,   readwrite); -- Bit15    Master Enable       (0=Disable, 1=Enable)
   
   constant SOUNDBIAS                                : regmap_type := (16#504#,   9,      0,        1, 16#0200#,   readwrite); -- (0..3FFh, usually 200h)

   constant SOUNDCAP                                 : regmap_type := (16#508#,  15,      0,        1,        0,   writeonly);
   constant SOUNDCAP0_Control                        : regmap_type := (16#508#,   0,      0,        1,        0,   readwrite); -- Bit0     Control of Associated Sound Channels (ANDed with Bit7) SNDCAP0CNT: Output Sound Channel 1 (0=As such, 1=Add to Channel 0) Caution: Addition mode works only if BOTH Bit0 and Bit7 are set.
   constant SOUNDCAP0_Capture_Source                 : regmap_type := (16#508#,   1,      1,        1,        0,   readwrite); -- Bit1     Capture Source Selection SNDCAP0CNT: Capture 0 Source (0=Left Mixer, 1=Channel 0/Bugged)
   constant SOUNDCAP0_Capture_Repeat                 : regmap_type := (16#508#,   2,      2,        1,        0,   readwrite); -- Bit2     Capture Repeat        (0=Loop, 1=One-shot)
   constant SOUNDCAP0_Capture_Format                 : regmap_type := (16#508#,   3,      3,        1,        0,   readwrite); -- Bit3     Capture Format        (0=PCM16, 1=PCM8)
   constant SOUNDCAP0_Capture_Start_Status           : regmap_type := (16#508#,   7,      7,        1,        0,   readwrite); -- Bit7     Capture Start/Status  (0=Stop, 1=Start/Busy)
   constant SOUNDCAP1_Control                        : regmap_type := (16#508#,   8,      8,        1,        0,   readwrite); -- Bit8     Control of Associated Sound Channels (ANDed with Bit7)  SNDCAP1CNT: Output Sound Channel 3 (0=As such, 1=Add to Channel 2) Caution: Addition mode works only if BOTH Bit0 and Bit7 are set.
   constant SOUNDCAP1_Capture_Source                 : regmap_type := (16#508#,   9,      9,        1,        0,   readwrite); -- Bit9     Capture Source Selection SNDCAP1CNT: Capture 1 Source (0=Right Mixer, 1=Channel 2/Bugged)
   constant SOUNDCAP1_Capture_Repeat                 : regmap_type := (16#508#,  10,     10,        1,        0,   readwrite); -- Bit10    Capture Repeat        (0=Loop, 1=One-shot)
   constant SOUNDCAP1_Capture_Format                 : regmap_type := (16#508#,  11,     11,        1,        0,   readwrite); -- Bit11    Capture Format        (0=PCM16, 1=PCM8)
   constant SOUNDCAP1_Capture_Start_Status           : regmap_type := (16#508#,  15,     15,        1,        0,   readwrite); -- Bit15    Capture Start/Status  (0=Stop, 1=Start/Busy)
   
   constant SNDCAP0DAD                               : regmap_type := (16#510#,  26,      0,        1,        0,   readwrite); -- Destination address (word aligned, bit0-1 are always zero)
   constant SNDCAP0LEN                               : regmap_type := (16#510#,  15,      0,        1,        0,   readwrite); -- Buffer length (1..FFFFh words) (ie. N*4 bytes)
   constant SNDCAP1DAD                               : regmap_type := (16#518#,  26,      0,        1,        0,   readwrite); -- Destination address (word aligned, bit0-1 are always zero)
   constant SNDCAP1LEN                               : regmap_type := (16#51C#,  15,      0,        1,        0,   readwrite); -- Buffer length (1..FFFFh words) (ie. N*4 bytes)


end package;